`ifndef SIPO_VH
`define SIPO_VH

`define MMIO_BASE_ADDR 32'h6000_0000
`define SIPO_DEPTH 256
`define SIPO_WIDTH 64
`define SYNC_STAGES 3

`endif /* SIPO_VH */
